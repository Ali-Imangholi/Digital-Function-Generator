`timescale 1ps/1ps
module AND(input in_and_1_ , input in_and_2_ , output out_and);
assign out_and  = and (in_and_1_ , in_and_2_);
endmodule